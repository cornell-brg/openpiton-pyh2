`timescale 1ns/1ps

module tbench_noc_axi4_bridge ;
wire m_axi_bready ;
wire m_axi_rready ;
wire m_axi_arvalid ;
wire [`AXI4_USER_WIDTH-1:0] m_axi_aruser ;
wire [`AXI4_REGION_WIDTH-1:0] m_axi_arregion ;
wire [`AXI4_QOS_WIDTH-1:0] m_axi_arqos ;
wire [`AXI4_PROT_WIDTH-1:0] m_axi_arprot ;
wire [`AXI4_CACHE_WIDTH-1:0] m_axi_arcache ;
wire m_axi_arlock ;
wire [`AXI4_BURST_WIDTH-1:0] m_axi_arburst ;
wire [`AXI4_SIZE_WIDTH-1:0] m_axi_arsize ;
wire [`AXI4_LEN_WIDTH-1:0] m_axi_arlen ;
wire [`AXI4_ADDR_WIDTH-1:0] m_axi_araddr ;
wire [`AXI4_ID_WIDTH-1:0] m_axi_arid ;
wire m_axi_wvalid ;
wire [`AXI4_USER_WIDTH-1:0] m_axi_wuser ;
wire m_axi_wlast ;
wire [`AXI4_STRB_WIDTH-1:0] m_axi_wstrb ;
wire [`AXI4_DATA_WIDTH-1:0] m_axi_wdata ;
wire [`AXI4_ID_WIDTH-1:0] m_axi_wid ;
wire m_axi_awvalid ;
wire [`AXI4_USER_WIDTH-1:0] m_axi_awuser ;
wire [`AXI4_REGION_WIDTH-1:0] m_axi_awregion ;
wire [`AXI4_QOS_WIDTH-1:0] m_axi_awqos ;
wire [`AXI4_PROT_WIDTH-1:0] m_axi_awprot ;
wire [`AXI4_CACHE_WIDTH-1:0] m_axi_awcache ;
wire m_axi_awlock ;
wire [`AXI4_BURST_WIDTH-1:0] m_axi_awburst ;
wire [`AXI4_SIZE_WIDTH-1:0] m_axi_awsize ;
wire [`AXI4_LEN_WIDTH-1:0] m_axi_awlen ;
wire [`AXI4_ADDR_WIDTH-1:0] m_axi_awaddr ;
wire [`AXI4_ID_WIDTH-1:0] m_axi_awid ;
wire [`NOC_DATA_WIDTH-1:0] bridge_dst_vr_noc3_dat ;
wire bridge_dst_vr_noc3_val ;
wire src_bridge_vr_noc2_rdy ;
reg m_axi_bvalid ;
reg [`AXI4_USER_WIDTH-1:0] m_axi_buser ;
reg [`AXI4_RESP_WIDTH-1:0] m_axi_bresp ;
reg [`AXI4_ID_WIDTH-1:0] m_axi_bid ;
reg m_axi_rvalid ;
reg [`AXI4_USER_WIDTH-1:0] m_axi_ruser ;
reg m_axi_rlast ;
reg [`AXI4_RESP_WIDTH-1:0] m_axi_rresp ;
reg [`AXI4_DATA_WIDTH-1:0] m_axi_rdata ;
reg [`AXI4_ID_WIDTH-1:0] m_axi_rid ;
reg m_axi_arready ;
reg m_axi_wready ;
reg m_axi_awready ;
reg bridge_dst_vr_noc3_rdy ;
reg [`NOC_DATA_WIDTH-1:0] src_bridge_vr_noc2_dat ;
reg src_bridge_vr_noc2_val ;
reg phy_init_done ;
reg uart_boot_en ;
reg reset ;
reg rst_n ;
reg clk ;
initial #9.852 $finish;
initial $dumpvars;
initial begin
    #0  m_axi_bvalid = 1'b0;
    #2.250  m_axi_bvalid = 1'b1;
    #0.100  m_axi_bvalid = 1'b0;
    #4.400  m_axi_bvalid = 1'b1;
    #0.100  m_axi_bvalid = 1'b0;
end
initial begin
    #0  m_axi_buser = 11'b00000000000;
end
initial begin
    #0  m_axi_bresp = 2'b00;
end
initial begin
    #0  m_axi_bid = 6'b000000;
    #6.750  m_axi_bid = 6'b000001;
    #0.100  m_axi_bid = 6'b000000;
end
initial begin
    #0  m_axi_rvalid = 1'b0;
    #2.450  m_axi_rvalid = 1'b1;
    #0.100  m_axi_rvalid = 1'b0;
    #0.500  m_axi_rvalid = 1'b1;
    #0.100  m_axi_rvalid = 1'b0;
    #0.200  m_axi_rvalid = 1'b1;
    #0.100  m_axi_rvalid = 1'b0;
    #0.500  m_axi_rvalid = 1'b1;
    #0.100  m_axi_rvalid = 1'b0;
    #0.900  m_axi_rvalid = 1'b1;
    #0.100  m_axi_rvalid = 1'b0;
    #0.900  m_axi_rvalid = 1'b1;
    #0.100  m_axi_rvalid = 1'b0;
end
initial begin
    #0  m_axi_ruser = 11'b00000000000;
end
initial begin
    #0  m_axi_rlast = 1'b0;
    #2.450  m_axi_rlast = 1'b1;
    #0.100  m_axi_rlast = 1'b0;
    #0.500  m_axi_rlast = 1'b1;
    #0.100  m_axi_rlast = 1'b0;
    #0.200  m_axi_rlast = 1'b1;
    #0.100  m_axi_rlast = 1'b0;
    #0.500  m_axi_rlast = 1'b1;
    #0.100  m_axi_rlast = 1'b0;
    #0.500  m_axi_rlast = 1'b1;
    #0.500  m_axi_rlast = 1'b0;
    #0.500  m_axi_rlast = 1'b1;
    #0.500  m_axi_rlast = 1'b0;
end
initial begin
    #0  m_axi_rresp = 2'b00;
end
initial begin
    #0  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    #2.450  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010110011101011000000001100;
    #0.100  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    #0.500  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010110011101011000000001100;
    #0.100  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    #0.200  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010110011101011000000001100;
    #0.100  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    #0.500  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010110011101011000000001100;
    #0.100  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    #0.500  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010110011101011000000001100;
    #0.500  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    #0.500  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010110011101011000000001100;
    #0.500  m_axi_rdata = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end
initial begin
    #0  m_axi_rid = 6'b000000;
    #2.450  m_axi_rid = 6'b000001;
    #0.100  m_axi_rid = 6'b000000;
    #0.800  m_axi_rid = 6'b000001;
    #0.100  m_axi_rid = 6'b000000;
    #1.100  m_axi_rid = 6'b000001;
    #0.500  m_axi_rid = 6'b000000;
end
initial begin
    #0  m_axi_arready = 1'b0;
    #0.250  m_axi_arready = 1'b1;
end
initial begin
    #0  m_axi_wready = 1'b0;
    #0.250  m_axi_wready = 1'b1;
end
initial begin
    #0  m_axi_awready = 1'b0;
    #0.250  m_axi_awready = 1'b1;
end
initial begin
    #0  bridge_dst_vr_noc3_rdy = 1'b0;
    #0.250  bridge_dst_vr_noc3_rdy = 1'b1;
end
initial begin
    #0  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    #0.250  src_bridge_vr_noc2_dat = 64'b0000000000001000000000000000000000000010100000111100000000000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000000010000000000000000011100000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000001000000010000000000000000000000000000000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000011111010110011101011000000001100;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    #0.700  src_bridge_vr_noc2_dat = 64'b0000000000001000000000000000000000000000100000111000000000000000;
    #0.200  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000000010000000000000000011100000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000001000000010000000000000000000000000000000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000001000000000000000000000000000100000111000000000000000;
    #0.200  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000000010000000000000000011100000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000001000000010000000000000000000000000000000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000001000000000000000000000000000100000111000000000000000;
    #0.200  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000000010000000000000000011100000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000001000000010000000000000000000000000000000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000001000000000000000000000000000100000111000000000000000;
    #0.200  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000000010000000000000000011100000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000001000000010000000000000000000000000000000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000001000000000000000000000000000100000111000000000000000;
    #0.200  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000000010000000000000000011100000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000001000000010000000000000000000000000000000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000001000000000000000000000000000100000111000000000000000;
    #0.200  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000000010000000000000000011100000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000001000000010000000000000000000000000000000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000001000000000000000000000000010100000111100000000000000;
    #0.200  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000000010000000000000000011100000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000001000000010000000000000000000000000000000000;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000010001011101011011111000000001101;
    #0.100  src_bridge_vr_noc2_dat = 64'b0000000000000000000000000000000000000000000000000000000000000000;
end
initial begin
    #0  src_bridge_vr_noc2_val = 1'b0;
    #0.250  src_bridge_vr_noc2_val = 1'b1;
    #1.100  src_bridge_vr_noc2_val = 1'b0;
    #0.100  src_bridge_vr_noc2_val = 1'b1;
    #0.300  src_bridge_vr_noc2_val = 1'b0;
    #0.100  src_bridge_vr_noc2_val = 1'b1;
    #0.300  src_bridge_vr_noc2_val = 1'b0;
    #0.100  src_bridge_vr_noc2_val = 1'b1;
    #0.300  src_bridge_vr_noc2_val = 1'b0;
    #0.100  src_bridge_vr_noc2_val = 1'b1;
    #0.300  src_bridge_vr_noc2_val = 1'b0;
    #0.100  src_bridge_vr_noc2_val = 1'b1;
    #0.300  src_bridge_vr_noc2_val = 1'b0;
    #0.100  src_bridge_vr_noc2_val = 1'b1;
    #0.300  src_bridge_vr_noc2_val = 1'b0;
    #0.100  src_bridge_vr_noc2_val = 1'b1;
    #1.100  src_bridge_vr_noc2_val = 1'b0;
end
initial begin
    #0  phy_init_done = 1'b0;
    #0.050  phy_init_done = 1'b1;
end
initial begin
    #0  uart_boot_en = 1'b0;
end
initial begin
    #0  reset = 1'b0;
    #0.050  reset = 1'b1;
    #0.200  reset = 1'b0;
end
initial begin
    #0  rst_n = 1'b0;
    #0.250  rst_n = 1'b1;
end
initial begin
     clk = 1'b0;
    forever #0.050  clk = ~ clk ;
end
noc_axi4_bridge noc_axi4_bridge (
    // Clock + Reset
    .clk( clk ),
    .rst_n( rst_n ),
    .reset( reset ),
    .uart_boot_en( uart_boot_en ),
    .phy_init_done( phy_init_done ),

    // Noc interface
    .src_bridge_vr_noc2_val( src_bridge_vr_noc2_val ),
    .src_bridge_vr_noc2_dat( src_bridge_vr_noc2_dat ),
    .src_bridge_vr_noc2_rdy( src_bridge_vr_noc2_rdy ),
    .bridge_dst_vr_noc3_val( bridge_dst_vr_noc3_val ),
    .bridge_dst_vr_noc3_dat( bridge_dst_vr_noc3_dat ),
    .bridge_dst_vr_noc3_rdy( bridge_dst_vr_noc3_rdy ),

    // AXI interface
    .m_axi_awid ( m_axi_awid ),
    .m_axi_awaddr ( m_axi_awaddr ),
    .m_axi_awlen ( m_axi_awlen ),
    .m_axi_awsize ( m_axi_awsize ),
    .m_axi_awburst ( m_axi_awburst ),
    .m_axi_awlock ( m_axi_awlock ),
    .m_axi_awcache ( m_axi_awcache ),
    .m_axi_awprot ( m_axi_awprot ),
    .m_axi_awqos ( m_axi_awqos ),
    .m_axi_awregion ( m_axi_awregion ),
    .m_axi_awuser ( m_axi_awuser ),
    .m_axi_awvalid ( m_axi_awvalid ),
    .m_axi_awready ( m_axi_awready ),

    .m_axi_wid( m_axi_wid ),
    .m_axi_wdata( m_axi_wdata ),
    .m_axi_wstrb( m_axi_wstrb ),
    .m_axi_wlast( m_axi_wlast ),
    .m_axi_wuser( m_axi_wuser ),
    .m_axi_wvalid( m_axi_wvalid ),
    .m_axi_wready( m_axi_wready ),

    .m_axi_arid( m_axi_arid ),
    .m_axi_araddr( m_axi_araddr ),
    .m_axi_arlen( m_axi_arlen ),
    .m_axi_arsize( m_axi_arsize ),
    .m_axi_arburst( m_axi_arburst ),
    .m_axi_arlock( m_axi_arlock ),
    .m_axi_arcache( m_axi_arcache ),
    .m_axi_arprot( m_axi_arprot ),
    .m_axi_arqos( m_axi_arqos ),
    .m_axi_arregion( m_axi_arregion ),
    .m_axi_aruser( m_axi_aruser ),
    .m_axi_arvalid( m_axi_arvalid ),
    .m_axi_arready( m_axi_arready ),

    .m_axi_rid( m_axi_rid ),
    .m_axi_rdata( m_axi_rdata ),
    .m_axi_rresp( m_axi_rresp ),
    .m_axi_rlast( m_axi_rlast ),
    .m_axi_ruser( m_axi_ruser ),
    .m_axi_rvalid( m_axi_rvalid ),
    .m_axi_rready( m_axi_rready ),

    .m_axi_bid( m_axi_bid ),
    .m_axi_bresp( m_axi_bresp ),
    .m_axi_buser( m_axi_buser ),
    .m_axi_bvalid( m_axi_bvalid ),
    .m_axi_bready( m_axi_bready )
);
endmodule
